 library ieee;
 use ieee.std_logic_1164.all;
 use ieee.std_logic_unsigned.all;
 
 entity div is
	generic( n1 : integer := 50000000;
		    n400 : integer := 12500);
	port( CLK : in std_logic;
		  Q1   : out std_logic;
		  Q400 : out std_logic);
end;

architecture bhv of div is
signal tempQ1 : std_logic;
signal tempQ400 : std_logic;
begin
	process(CLK)
	variable num : integer range 0 to n1;
	begin
		if( rising_edge(CLK) ) then
			num := num + 1;
		end if;
		if( num <= n1/2 ) then
			tempQ1 <= '0';
		else
			tempQ1 <= '1';
		end if;
		if( num > n1 ) then	--清零
			num := 0;
		end if;
	end process;
	
	process(CLK)
	variable num : integer range 0 to n400;
	begin
		if( rising_edge(CLK) ) then
			num := num + 1;
		end if;
		if( num <= n400/2 ) then
			tempQ400 <= '0';
		else
			tempQ400 <= '1';
		end if;
		if( num > n400 ) then
			num := 0;
		end if;
	end process;
	Q1 <= tempQ1;
	Q400 <= tempQ400;
end architecture;